----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/18/2017 12:51:13 PM
-- Design Name: 
-- Module Name: reg - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity reg is
  Port (      D : in std_logic_vector(7 downto 0);
         CLK,LD : in std_logic;
              Q : out std_logic_vector(7 downto 0));
end reg;

architecture Behavioral of reg is

begin
    process (D, CLK, LD)
    begin
        if (rising_edge(CLK)) then
            if(LD = '1') then
                Q <= D;
            end if;
         end if;
      end process;

end Behavioral;
